 library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity prom_DMH is
    port (
		S: in STD_LOGIC_VECTOR (7 downto 0);
		clr: in std_logic;
        addr: in STD_LOGIC_VECTOR (7 downto 0);
        M: out STD_LOGIC_VECTOR (0 to 38)
    );
end prom_DMH;

architecture prom_DMH of prom_DMH is
type rom_array is array (NATURAL range <>) of STD_LOGIC_VECTOR (0 to 38);
type rom1_array is array (NATURAL range <>) of STD_LOGIC_VECTOR (0 to 38);
type rom2_array is array (NATURAL range <>) of STD_LOGIC_VECTOR (0 to 38);
type rom3_array is array (NATURAL range <>) of STD_LOGIC_VECTOR (0 to 38);
type rom4_array is array (NATURAL range <>) of STD_LOGIC_VECTOR (0 to 38);
type rom5_array is array (NATURAL range <>) of STD_LOGIC_VECTOR (0 to 38);
type rom6_array is array (NATURAL range <>) of STD_LOGIC_VECTOR (0 to 38);
type rom7_array is array (NATURAL range <>) of STD_LOGIC_VECTOR (0 to 38);
type rom8_array is array (NATURAL range <>) of STD_LOGIC_VECTOR (0 to 38);
type rom9_array is array (NATURAL range <>) of STD_LOGIC_VECTOR (0 to 38);
type rom10_array is array (NATURAL range <>) of STD_LOGIC_VECTOR (0 to 38);
type rom11_array is array (NATURAL range <>) of STD_LOGIC_VECTOR (0 to 38);
type rom12_array is array (NATURAL range <>) of STD_LOGIC_VECTOR (0 to 38);
type rom13_array is array (NATURAL range <>) of STD_LOGIC_VECTOR (0 to 38);
type rom14_array is array (NATURAL range <>) of STD_LOGIC_VECTOR (0 to 38);
type rom15_array is array (NATURAL range <>) of STD_LOGIC_VECTOR (0 to 38);
type rom16_array is array (NATURAL range <>) of STD_LOGIC_VECTOR (0 to 38);
type rom17_array is array (NATURAL range <>) of STD_LOGIC_VECTOR (0 to 38);
type rom18_array is array (NATURAL range <>) of STD_LOGIC_VECTOR (0 to 38);
type rom19_array is array (NATURAL range <>) of STD_LOGIC_VECTOR (0 to 38);
type rom20_array is array (NATURAL range <>) of STD_LOGIC_VECTOR (0 to 38);
type rom21_array is array (NATURAL range <>) of STD_LOGIC_VECTOR (0 to 38);
type rom22_array is array (NATURAL range <>) of STD_LOGIC_VECTOR (0 to 38);
type rom23_array is array (NATURAL range <>) of STD_LOGIC_VECTOR (0 to 38);	
type rom24_array is array (NATURAL range <>) of STD_LOGIC_VECTOR (0 to 38);

constant rom: rom_array := (
	"000000000000000000000000000000000000000",		--0
	"000000000000000000000000000000000000000",		--1
	"000000000000000000010000000000000000000", 		--2
	"000000000000000000101000000000000000000", 		--3
	"000000000000000001000100000000000000000", 		--4
	"000000000000000010000010000000000000000", 		--5
	"000000000000000100000001000000000000000", 		--6
	"000000000000001000000000100000000000000", 		--7
	"000000000000010000000000010000000000000", 		--8
	"000000000000100000000000001000000000000", 		--9
	"000000000001000000000000000100000000000", 		--10
	"000000000010000000000000000010000000000", 		--11
	"000000000100000000000000000001000000000", 		--12
	"000000001000000000000000000000100000000", 		--13
	"000000011111111111111111111111110000000", 		--14
	"000000100000000000000000000000001000000", 		--15
	"000001000000000000000000000000000100000", 		--16
	"000010000000000000000000000000000010000",	 	--17 
	"000000000000000000000000000000000000000",		--18
	"000000000000000000000000000000000000000",		--19
	"000000000000000000000000000000000000000"		--20
	);

constant rom1: rom1_array := (
	"000000000000000000000000000000000000000",		--0
	"000000000000000000000000000000000000000",		--1
	"000000000000000000000000000000000000000", 		--2
	"000000000000000011100000000000000000000", 		--3
	"000000000000000010110000000000000000000", 		--4
	"000000000000001100011000000000000000000", 		--5
	"000000000000001000000100000000000000000", 		--6
	"000000000000011000000011000000000000000", 		--7
	"000000000000110000000001100000000000000", 		--8
	"000000000001100000000000011000000000000", 		--9
	"000000000001100000000000001100000000000", 		--10
	"000000000011000000000000000110000000000", 		--11
	"000000000010000000000000000001100000000", 		--12
	"000000000100000000000000000000110000000", 		--13
	"000000001000000000011111111111111000000", 		--14
	"000000011111111111111000000000001100000", 		--15
	"000000010000000000000000000000000011000", 		--16
	"000000110000000000000000000000000001000",	 	--17 
	"000001100000000000000000000000000000000",	   	--18
	"000000000000000000000000000000000000000",		--19
	"000000000000000000000000000000000000000"		--20
	);

constant rom2: rom2_array := ( 
	"000000000000000000000000000000000000000",		--0
	"000000000000000000000000000000000000000",		--1
	"000000000000000000000000000000000000000", 		--2
	"000000000000001110000000000000000000000", 		--3
	"000000000000001101100000000000000000000", 		--4
	"000000000000001000110000000000000000000", 		--5
	"000000000000010000001100000000000000000", 		--6
	"000000000000010000000011000000000000000", 		--7
	"000000000000110000000001100000000000000", 		--8
	"000000000001100000000000011000000000000", 		--9
	"000000000001100000000000000110000000000", 		--10
	"000000000011000000000000000001100000000", 		--11
	"000000000010000000000000000000110000000", 		--12
	"000000000110000000000000000001111000000", 		--13
	"000000000100000000011111111111111100000", 		--14
	"000000001111111111111000000000000011000", 		--15
	"000000001000000000000000000000000001000", 		--16
	"000000011000000000000000000000000000000",	 	--17 
	"000000010000000000000000000000000000000",		--18
	"000000110000000000000000000000000000000",		--19
	"000000000000000000000000000000000000000"		--20
	);

constant rom3: rom3_array := (
	"000000000000000000000000000000000000000",		--0
	"000000000000000000000000000000000000000",		--1
	"000000000000000000000000000000000000000", 		--2
	"000000000000110000000000000000000000000", 		--3
	"000000000000110110000000000000000000000", 		--4
	"000000000000110011100000000000000000000", 		--5
	"000000000000100000110000000000000000000", 		--6
	"000000000000100000001110000000000000000", 		--7
	"000000000001100000000011100000000000000", 		--8
	"000000000001100000000000111000000000000", 		--9
	"000000000001000000000000000110000000000", 		--10
	"000000000011000000000000000001100000000", 		--11
	"000000000011000000000000000000111000000", 		--12
	"000000000010000000000000001111111110000", 		--13
	"000000000010000000011111111110000011000", 		--14
	"000000000111111111110000000000000000110", 		--15
	"000000000111100000000000000000000000000", 		--16
	"000000000100000000000000000000000000000",	 	--17 
	"000000000100000000000000000000000000000",		--18
	"000000001100000000000000000000000000000",		--19
	"000000000000000000000000000000000000000"		--20
	);

constant rom4: rom4_array := (
	"000000000000000000000000000000000000000",		--0
	"000000000000000000000000000000000000000",		--1
	"000000000000000000000000000000000000000", 		--2
	"000000000011000000000000000000000000000", 		--3
	"000000000011110000000000000000000000000", 		--4
	"000000000011001110000000000000000000000", 		--5
	"000000000011000001110000000000000000000", 		--6
	"000000000011000000001100000000000000000", 		--7
	"000000000010000000000011000000000000000", 		--8
	"000000000010000000000000011000000000000", 		--9
	"000000000010000000000000000111000000000", 		--10
	"000000000010000000000000000001110000000", 		--11
	"000000000010000000000000000011111100000", 		--12
	"000000000010000000000000111111000011100", 		--13
	"000000000010000000111111100000000000110", 		--14
	"000000000110111111110000000000000000000", 		--15
	"000000000111111000000000000000000000000", 		--16
	"000000000110000000000000000000000000000",	 	--17 
	"000000000110000000000000000000000000000",		--18
	"000000000110000000000000000000000000000",		--19
	"000000000100000000000000000000000000000"		--20
	);

constant rom5: rom5_array := (
	"000000000000000000000000000000000000000",		--0
	"000000000000000000000000000000000000000",		--1
	"000000000000000000000000000000000000000", 		--2
	"000000001100000000000000000000000000000", 		--3
	"000000001111100000000000000000000000000", 		--4
	"000000001100011100000000000000000000000", 		--5
	"000000000100000011100000000000000000000", 		--6
	"000000000110000000011110000000000000000", 		--7
	"000000000110000000000001110000000000000", 		--8
	"000000000110000000000000001111000000000", 		--9
	"000000000010000000000000000001110000000", 		--10
	"000000000010000000000000000011111110000", 		--11
	"000000000010000000000000011111000001110", 		--12
	"000000000011000000000111110000000000001", 		--13
	"000000000011000000111100000000000000000", 		--14
	"000000000001011111110000000000000000000", 		--15
	"000000000001111000000000000000000000000", 		--16
	"000000000001100000000000000000000000000",	 	--17 
	"000000000001100000000000000000000000000",		--18
	"000000000001100000000000000000000000000",		--19
	"000000000001100000000000000000000000000"		--20
	);

constant rom6: rom6_array := (
	"000000000000000000000000000000000000000",		--0
	"000000000000000000000000000000000000000",		--1
	"000000000000000000000000000000000000000", 		--2
	"000000000000000000000000000000000000000", 		--3
	"000000111100000000000000000000000000000", 		--4
	"000000110011110000000000000000000000000", 		--5
	"000000010000001111000000000000000000000", 		--6
	"000000011000000000011110000000000000000", 		--7
	"000000001000000000000001110000000000000", 		--8
	"000000001100000000000000001111000000000", 		--9
	"000000000100000000000000000001111100000", 		--10
	"000000000010000000000000001111100011110", 		--11
	"000000000010000000000000111100000000010", 		--12
	"000000000011000000001111100000000000000", 		--13
	"000000000011000001111100000000000000000", 		--14
	"000000000001001111100000000000000000000", 		--15
	"000000000001111000000000000000000000000", 		--16
	"000000000000100000000000000000000000000",	 	--17 
	"000000000000110000000000000000000000000",		--18
	"000000000000110000000000000000000000000",		--19
	"000000000000010000000000000000000000000"		--20
	);

constant rom7: rom7_array := (	
	"000000000000000000000000000000000000000",		--0
	"000000000000000000000000000000000000000",		--1
	"000000000000000000000000000000000000000", 		--2
	"000000000000000000000000000000000000000", 		--3
	"000000000000000000000000000000000000000", 		--4
	"000011111110000000000000000000000000000", 		--5
	"000001100001111110000000000000000000000", 		--6
	"000000100000000001111110000000000000000", 		--7
	"000000010000000000000001111110000000000", 		--8
	"000000001000000000000000000001111110000", 		--9
	"000000001100000000000000000111100001110", 		--10
	"000000000110000000000000011110000000000", 		--11
	"000000000010000000000001110000000000000", 		--12
	"000000000011000000001111000000000000000", 		--13
	"000000000001100000111100000000000000000", 		--14
	"000000000000110011110000000000000000000", 		--15
	"000000000000111111000000000000000000000", 		--16
	"000000000000011100000000000000000000000",	 	--17 
	"000000000000001100000000000000000000000",		--18
	"000000000000000110000000000000000000000",		--19
	"000000000000000010000000000000000000000"		--20
	);

constant rom8: rom8_array := ( 
	"000000000000000000000000000000000000000",		--0
	"000000000000000000000000000000000000000",		--1
	"000000000000000000000000000000000000000", 		--2
	"000000000000000000000000000000000000000", 		--3
	"000000000000000000000000000000000000000", 		--4
	"001110000000000000000000000000000000000", 		--5
	"000110111111111000000000000000000000000", 		--6
	"000011000000000111111111111000000000000", 		--7
	"000001100000000000000000001111111111000", 		--8
	"000000110000000000000000000111100001110", 		--9
	"000000011000000000000000001110000000000", 		--10
	"000000001100000000000000111000000000000", 		--11
	"000000000110000000000011110000000000000", 		--12
	"000000000001100000001111000000000000000", 		--13
	"000000000000110000011110000000000000000", 		--14
	"000000000000011001111000000000000000000", 		--15
	"000000000000011111100000000000000000000", 		--16
	"000000000000000110000000000000000000000",	 	--17 
	"000000000000000011000000000000000000000",		--18
	"000000000000000001100000000000000000000",		--19
	"000000000000000000110000000000000000000"		--20
	);

constant rom9: rom9_array := (
	"000000000000000000000000000000000000000",		--0
	"000000000000000000000000000000000000000",		--1
	"000000000000000000000000000000000000000", 		--2
	"000000000000000000000000000000000000000", 		--3
	"000000000000000000000000000000000000000", 		--4
	"000000000000000000000000000000000000000", 		--5
	"011111111111111111110000000000000000000", 		--6
	"001100000000000000011111111111111111100", 		--7
	"000011000000000000000000000111000000000", 		--8
	"000001100000000000000000001110000000000", 		--9
	"000000011000000000000000011100000000000", 		--10
	"000000001100000000000001111000000000000", 		--11
	"000000000111000000000011100000000000000", 		--12
	"000000000001100000001111000000000000000", 		--13
	"000000000000011000011110000000000000000", 		--14
	"000000000000001100111000000000000000000", 		--15
	"000000000000000111110000000000000000000", 		--16
	"000000000000000001100000000000000000000",	 	--17 
	"000000000000000000110000000000000000000",		--18
	"000000000000000000001100000000000000000",		--19
	"000000000000000000000100000000000000000"		--20
	);

constant rom10: rom10_array := ( 
	"000000000000000000000000000000000000000",		--0
	"000000000000000000000000000000000000000",		--1
	"000000000000000000000000000000000000000", 		--2
	"000000000000000000000000000000000000000", 		--3
	"000000000000000000000000000000000000000", 		--4
	"000000000000000000000000000000000000000", 		--5
	"000000000000000011111111111111111111100", 		--6
	"111111111111111100000000000111000000000", 		--7
	"001100000000000000000000001110000000000", 		--8
	"000011000000000000000000011100000000000", 		--9
	"000000110000000000000000011100000000000", 		--10
	"000000001100000000000000111000000000000", 		--11
	"000000000111000000000001100000000000000", 		--12
	"000000000000110000000011100000000000000", 		--13
	"000000000000001110000111000000000000000", 		--14
	"000000000000000011101110000000000000000", 		--15
	"000000000000000000111100000000000000000", 		--16
	"000000000000000000001110000000000000000",	 	--17 
	"000000000000000000000011100000000000000",		--18
	"000000000000000000000000110000000000000",		--19
	"000000000000000000000000000000000000000"		--20
	);

constant rom11: rom11_array := ( 
	"000000000000000000000000000000000000000",		--0
	"000000000000000000000000000000000000000",		--1
	"000000000000000000000000000000000000000", 		--2
	"000000000000000000000000000000000000000", 		--3
	"000000000000000000000000000000011111000", 		--4
	"000000000000000000000001111111110000000", 		--5
	"000000000000000000111111000110000000000", 		--6
	"000000000000111111000000001110000000000", 		--7
	"000000111111000000000000001110000000000", 		--8
	"011111000000000000000000001100000000000", 		--9
	"001111000000000000000000011100000000000", 		--10
	"000000111000000000000000011100000000000", 		--11
	"000000000111100000000000011000000000000", 		--12
	"000000000000111000000000011000000000000", 		--13
	"000000000000000011110000111000000000000", 		--14
	"000000000000000000011110111000000000000", 		--15
	"000000000000000000000001110000000000000", 		--16
	"000000000000000000000000001111000000000",	 	--17 
	"000000000000000000000000000001110000000",		--18
	"000000000000000000000000000000000000000",		--19
	"000000000000000000000000000000000000000"		--20
	);

constant rom12: rom12_array := (
	"000000000000000000000000000000000000000",		--0
	"000000000000000000000000000000000000000",		--1
	"000000000000000000000000000000000000000", 		--2
	"000000000000000000000000000000011110000", 		--3
	"000000000000000000000000000111110000000", 		--4
	"000000000000000000000111111110000000000", 		--5
	"000000000000000000111110001110000000000", 		--6
	"000000000000001111000000001100000000000", 		--7
	"000000000111100000000000001100000000000", 		--8
	"000011111000000000000000001100000000000", 		--9
	"001110000000000000000000001100000000000", 		--10
	"000111110000000000000000001100000000000", 		--11
	"000000001111000000000000001100000000000", 		--12
	"000000000000111110000000001100000000000", 		--13
	"000000000000000001111000001100000000000", 		--14
	"000000000000000000000111101100000000000", 		--15
	"000000000000000000000000011111100000000", 		--16
	"000000000000000000000000000000111100000",	 	--17 
	"000000000000000000000000000000000000000",		--18
	"000000000000000000000000000000000000000",		--19
	"000000000000000000000000000000000000000"		--20
	);
constant rom13: rom13_array := (
	"000000000000000000000000000000000000000", 		--0
	"000000000000000000000000000000000000000", 		--1
	"000000000000000000000000000001110000000", 		--2
	"000000000000000000000000001111000000000", 		--3
	"000000000000000000000001110000000000000", 		--4
	"000000000000000000011110111000000000000", 		--5
	"000000000000000011110000111000000000000", 		--6
	"000000000000111000000000011000000000000", 		--7
	"000000000111100000000000011000000000000", 		--8
	"000000111000000000000000011100000000000", 		--9
	"001111000000000000000000011100000000000", 		--10
	"011111000000000000000000001100000000000", 		--11
	"000000111111000000000000001110000000000", 		--12
	"000000000000111111000000001110000000000", 		--13
	"000000000000000000111111000110000000000", 		--14
	"000000000000000000000001111111110000000",	 	--15 
	"000000000000000000000000000000011111000",		--16
	"000000000000000000000000000000000000000",		--17
	"000000000000000000000000000000000000000",		--18
	"000000000000000000000000000000000000000",		--19
	"000000000000000000000000000000000000000"		--20
	); 
constant rom14: rom14_array := (
	"000000000000000000000000000000000000000",		--0
	"000000000000000000000000110000000000000",		--1
	"000000000000000000000011100000000000000", 		--2
	"000000000000000000001110000000000000000", 		--3
	"000000000000000000111100000000000000000", 		--4
	"000000000000000011101110000000000000000", 		--5
	"000000000000001110000111000000000000000", 		--6
	"000000000000110000000011100000000000000", 		--7
	"000000000111000000000001100000000000000", 		--8
	"000000001100000000000000111000000000000", 		--9
	"000000110000000000000000011100000000000", 		--10
	"000011000000000000000000011100000000000", 		--11
	"001100000000000000000000001110000000000", 		--12
	"111111111111111100000000000111000000000", 		--13
	"000000000000000011111111111111111111100", 		--14
	"000000000000000000000000000000000000000", 		--15
	"000000000000000000000000000000000000000", 		--16
	"000000000000000000000000000000000000000",	 	--17 
	"000000000000000000000000000000000000000",		--18
	"000000000000000000000000000000000000000",		--19
	"000000000000000000000000000000000000000"		--20
	);
constant rom15: rom15_array := (
	"000000000000000000000100000000000000000",		--0
	"000000000000000000001100000000000000000",		--1
	"000000000000000000110000000000000000000", 		--2
	"000000000000000001100000000000000000000", 		--3
	"000000000000000111110000000000000000000", 		--4
	"000000000000001100111000000000000000000", 		--5
	"000000000000011000011110000000000000000", 		--6
	"000000000001100000001111000000000000000", 		--7
	"000000000111000000000011100000000000000", 		--8
	"000000001100000000000001111000000000000", 		--9
	"000000011000000000000000011100000000000", 		--10
	"000001100000000000000000001110000000000", 		--11
	"000011000000000000000000000111000000000", 		--12
	"001100000000000000011111111111111111100", 		--13
	"011111111111111111110000000000000000000", 		--14
	"000000000000000000000000000000000000000", 		--15
	"000000000000000000000000000000000000000", 		--16
	"000000000000000000000000000000000000000",	 	--17 
	"000000000000000000000000000000000000000",		--18
	"000000000000000000000000000000000000000",		--19
	"000000000000000000000000000000000000000"		--20
	);
constant rom16: rom16_array := (
	"000000000000000000110000000000000000000",		--0
	"000000000000000001100000000000000000000",		--1
	"000000000000000011000000000000000000000", 		--2
	"000000000000000110000000000000000000000", 		--3
	"000000000000011111100000000000000000000", 		--4
	"000000000000011001111000000000000000000", 		--5
	"000000000000110000011110000000000000000", 		--6
	"000000000001100000001111000000000000000", 		--7
	"000000000110000000000011110000000000000", 		--8
	"000000001100000000000000111000000000000", 		--9
	"000000011000000000000000001110000000000", 		--10
	"000000110000000000000000000111100001110", 		--11
	"000001100000000000000000001111111111000", 		--12
	"000011000000000111111111111000000000000", 		--13
	"000110111111111000000000000000000000000", 		--14
	"001110000000000000000000000000000000000", 		--15
	"000000000000000000000000000000000000000", 		--16
	"000000000000000000000000000000000000000",	 	--17 
	"000000000000000000000000000000000000000",		--18
	"000000000000000000000000000000000000000",		--19
	"000000000000000000000000000000000000000"		--20
	);
constant rom17: rom17_array := (
	"000000000000000010000000000000000000000",		--0
	"000000000000000110000000000000000000000",		--1
	"000000000000001100000000000000000000000", 		--2
	"000000000000011100000000000000000000000", 		--3
	"000000000000111111000000000000000000000", 		--4
	"000000000000110011110000000000000000000", 		--5
	"000000000001100000111100000000000000000", 		--6
	"000000000011000000001111000000000000000", 		--7
	"000000000010000000000001110000000000000", 		--8
	"000000000110000000000000011110000000000", 		--9
	"000000001100000000000000000111100001110", 		--10
	"000000001000000000000000000001111110000", 		--11
	"000000010000000000000001111110000000000", 		--12
	"000000100000000001111110000000000000000", 		--13
	"000001100001111110000000000000000000000", 		--14
	"000011111110000000000000000000000000000", 		--15
	"000000000000000000000000000000000000000", 		--16
	"000000000000000000000000000000000000000",	 	--17 
	"000000000000000000000000000000000000000",		--18
	"000000000000000000000000000000000000000",		--19
	"000000000000000000000000000000000000000"		--20
	);
constant rom18: rom18_array := (
	"000000000000010000000000000000000000000",		--0
	"000000000000110000000000000000000000000",		--1
	"000000000000110000000000000000000000000", 		--2
	"000000000000100000000000000000000000000", 		--3
	"000000000001111000000000000000000000000", 		--4
	"000000000001001111100000000000000000000", 		--5
	"000000000011000001111100000000000000000", 		--6
	"000000000011000000001111100000000000000", 		--7
	"000000000010000000000000111100000000010", 		--8
	"000000000010000000000000001111100011110", 		--9
	"000000000100000000000000000001111100000", 		--10
	"000000001100000000000000001111000000000", 		--11
	"000000001000000000000001110000000000000", 		--12
	"000000011000000000011110000000000000000", 		--13
	"000000010000001111000000000000000000000", 		--14
	"000000110011110000000000000000000000000", 		--15
	"000000111100000000000000000000000000000", 		--16
	"000000000000000000000000000000000000000",	 	--17 
	"000000000000000000000000000000000000000",		--18
	"000000000000000000000000000000000000000",		--19
	"000000000000000000000000000000000000000"		--20
	);
constant rom19: rom19_array := (
	"000000000001100000000000000000000000000",		--0
	"000000000001100000000000000000000000000",		--1
	"000000000001100000000000000000000000000", 		--2
	"000000000001100000000000000000000000000", 		--3
	"000000000001111000000000000000000000000", 		--4
	"000000000001011111110000000000000000000", 		--5
	"000000000011000000111100000000000000000", 		--6
	"000000000011000000000111110000000000001", 		--7
	"000000000010000000000000011111000001110", 		--8
	"000000000010000000000000000011111110000", 		--9
	"000000000010000000000000000001110000000", 		--10
	"000000000110000000000000001111000000000", 		--11
	"000000000110000000000001110000000000000", 		--12
	"000000000110000000011110000000000000000", 		--13
	"000000000100000011100000000000000000000", 		--14
	"000000001100011100000000000000000000000", 		--15
	"000000001111100000000000000000000000000", 		--16
	"000000001100000000000000000000000000000",	 	--17 
	"000000000000000000000000000000000000000",		--18
	"000000000000000000000000000000000000000",		--19
	"000000000000000000000000000000000000000"		--20
	);
constant rom20: rom20_array := (
	"000000000100000000000000000000000000000",		--0
	"000000000110000000000000000000000000000",		--1
	"000000000110000000000000000000000000000", 		--2
	"000000000110000000000000000000000000000", 		--3
	"000000000111111000000000000000000000000", 		--4
	"000000000110111111110000000000000000000", 		--5
	"000000000010000000111111100000000000110", 		--6
	"000000000010000000000000111111000011100", 		--7
	"000000000010000000000000000011111100000", 		--8
	"000000000010000000000000000001110000000", 		--9
	"000000000010000000000000000111000000000", 		--10
	"000000000010000000000000011000000000000", 		--11
	"000000000010000000000011000000000000000", 		--12
	"000000000011000000001100000000000000000", 		--13
	"000000000011000001110000000000000000000", 		--14
	"000000000011001110000000000000000000000", 		--15
	"000000000011110000000000000000000000000", 		--16
	"000000000011000000000000000000000000000",	 	--17 
	"000000000000000000000000000000000000000",		--18
	"000000000000000000000000000000000000000",		--19
	"000000000000000000000000000000000000000"		--20
	);
constant rom21: rom21_array := (
	"000000000000000000000000000000000000000",		--0
	"000000001100000000000000000000000000000",		--1
	"000000000100000000000000000000000000000", 		--2
	"000000000100000000000000000000000000000", 		--3
	"000000000111100000000000000000000000000", 		--4
	"000000000111111111110000000000000000110", 		--5
	"000000000010000000011111111110000011000", 		--6
	"000000000010000000000000001111111110000", 		--7
	"000000000011000000000000000000111000000", 		--8
	"000000000011000000000000000001100000000", 		--9
	"000000000001000000000000000110000000000", 		--10
	"000000000001100000000000111000000000000", 		--11
	"000000000001100000000011100000000000000", 		--12
	"000000000000100000001110000000000000000", 		--13
	"000000000000100000110000000000000000000", 		--14
	"000000000000110011100000000000000000000", 		--15
	"000000000000110110000000000000000000000", 		--16
	"000000000000110000000000000000000000000",	 	--17 
	"000000000000000000000000000000000000000",		--18
	"000000000000000000000000000000000000000",		--19
	"000000000000000000000000000000000000000"		--20
	);
constant rom22: rom22_array := (
	"000000000000000000000000000000000000000",		--0
	"000000110000000000000000000000000000000",		--1
	"000000010000000000000000000000000000000", 		--2
	"000000011000000000000000000000000000000", 		--3
	"000000001000000000000000000000000001000", 		--4
	"000000001111111111111000000000000011000", 		--5
	"000000000100000000011111111111111100000", 		--6
	"000000000110000000000000000001111000000", 		--7
	"000000000010000000000000000000110000000", 		--8
	"000000000011000000000000000001100000000", 		--9
	"000000000001100000000000000110000000000", 		--10
	"000000000001100000000000011000000000000", 		--11
	"000000000000110000000001100000000000000", 		--12
	"000000000000010000000011000000000000000", 		--13
	"000000000000010000001100000000000000000", 		--14
	"000000000000001000110000000000000000000", 		--15
	"000000000000001101100000000000000000000", 		--16
	"000000000000001110000000000000000000000",	 	--17 
	"000000000000000000000000000000000000000",		--18
	"000000000000000000000000000000000000000",		--19
	"000000000000000000000000000000000000000"		--20
	); 
constant rom23: rom23_array := (
	"000000000000000000000000000000000000000",		--0
	"000000000000000000000000000000000000000",		--1
	"000001100000000000000000000000000000000", 		--2
	"000000110000000000000000000000000001000", 		--3
	"000000010000000000000000000000000011000", 		--4
	"000000011111111111111000000000001100000", 		--5
	"000000001000000000011111111111111000000", 		--6
	"000000000100000000000000000000110000000", 		--7
	"000000000010000000000000000001100000000", 		--8
	"000000000011000000000000000110000000000", 		--9
	"000000000001100000000000001100000000000", 		--10
	"000000000001100000000000011000000000000", 		--11
	"000000000000110000000001100000000000000", 		--12
	"000000000000011000000011000000000000000", 		--13
	"000000000000001000000100000000000000000", 		--14
	"000000000000001100011000000000000000000", 		--15
	"000000000000000010110000000000000000000", 		--16
	"000000000000000011100000000000000000000",	 	--17 
	"000000000000000000000000000000000000000",		--18
	"000000000000000000000000000000000000000",		--19
	"000000000000000000000000000000000000000"		--20
	);
constant rom24: rom24_array := (
	"000000000000000000000000000000000000000",		--0
	"000000000000000000000000000000000000000",		--1
	"000000000000000000000000000000000000000", 		--2
	"000010000000000000000000000000000010000", 		--3
	"000001000000000000000000000000000100000", 		--4
	"000000100000000000000000000000001000000", 		--5
	"000000011111111111111111111111110000000", 		--6
	"000000001000000000000000000000100000000", 		--7
	"000000000100000000000000000001000000000", 		--8
	"000000000010000000000000000010000000000", 		--9
	"000000000001000000000000000100000000000", 		--10
	"000000000000100000000000001000000000000", 		--11
	"000000000000010000000000010000000000000", 		--12
	"000000000000001000000000100000000000000", 		--13
	"000000000000000100000001000000000000000", 		--14
	"000000000000000010000010000000000000000", 		--15
	"000000000000000001000100000000000000000", 		--16
	"000000000000000000101000000000000000000",	 	--17 
	"000000000000000000010000000000000000000",		--18
	"000000000000000000000000000000000000000",		--19
	"000000000000000000000000000000000000000"		--20
	);
begin
	process(S,addr,clr)
	variable j: integer;
	begin 
		if clr = '1' then
    	 j := conv_integer(addr);
   		 M <= rom(j);
		elsif s = "00000000" then
		 j := conv_integer(addr);
   		 M <= rom(j);
		elsif s = "00000001" then
		 j := conv_integer(addr);
   		 M <= rom1(j);
		elsif s = "00000010" then
		 j := conv_integer(addr);
   		 M <= rom2(j);
		elsif s = "00000011" then
		 j := conv_integer(addr);
   		 M <= rom3(j);			
		elsif s = "00000100" then
		 j := conv_integer(addr);
   		 M <= rom4(j);			
		elsif s = "00000101" then
		 j := conv_integer(addr);
   		 M <= rom5(j);
		elsif s = "00000110" then
		 j := conv_integer(addr);
   		 M <= rom6(j);			
		elsif s = "00000111" then
		 j := conv_integer(addr);
   		 M <= rom7(j);			 
		elsif s = "00001000" then
		 j := conv_integer(addr);
   		 M <= rom8(j);			
		elsif s = "00001001" then
		 j := conv_integer(addr);
   		 M <= rom9(j);			
		elsif s = "00001010" then
		 j := conv_integer(addr);
   		 M <= rom10(j);			
		elsif s = "00001011" then
		 j := conv_integer(addr);
   		 M <= rom11(j);			
		elsif s = "00001100" then
		 j := conv_integer(addr);
   		 M <= rom12(j);	
		elsif s = "00001101" then
		 j := conv_integer(addr);
   		 M <= rom13(j);
		elsif s = "00001110" then
		 j := conv_integer(addr);
   		 M <= rom14(j);	
		elsif s = "00001111" then
		 j := conv_integer(addr);
   		 M <= rom15(j);	
		elsif s = "00010000" then
		 j := conv_integer(addr);
   		 M <= rom16(j);	
		elsif s = "00010001" then
		 j := conv_integer(addr);
   		 M <= rom17(j);	
		elsif s = "00010010" then
		 j := conv_integer(addr);
   		 M <= rom18(j);	
		elsif s = "00010011" then
		 j := conv_integer(addr);
   		 M <= rom19(j);	
		elsif s = "00010100" then
		 j := conv_integer(addr);
   		 M <= rom20(j);	
		elsif s = "00010101" then
		 j := conv_integer(addr);
   		 M <= rom21(j);	
		elsif s = "00010110" then
		 j := conv_integer(addr);
   		 M <= rom22(j);	
		elsif s = "00010111" then
		 j := conv_integer(addr);
   		 M <= rom23(j);	
		elsif s = "00011000" then
		 j := conv_integer(addr);
   		 M <= rom24(j);	
		end if;	
			
  end process;

end prom_DMH;