 library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity prom2_asteroid is
    port ( 

		rom_addra  : in std_logic_vector(7 downto 0);
        D: out STD_LOGIC_VECTOR (0 to 60)
    );
end prom2_asteroid;

architecture prom2_asteroid of prom2_asteroid is   
type rom_array is array (NATURAL range <>) of STD_LOGIC_VECTOR (0 to 60);
constant rom: rom_array := (   
	"0000000000000000000000001111111111111000000000000000000000000",		--0
	"0000000000000000000000110000000000000110000000000000000000000",		--1
	"0000000000000000000011000000000000000001111111110000000000000", 		--2
	"0000000000000000001100000000000000000000000000001110000000000", 		--3
	"0000000000000000110000000000000000000000000000000001100000000", 		--4
	"0000000000000111000000000000000000000000000000000000010000000", 		--5
	"0000000000111000000000000000000000000000000000000000010000000", 		--6
	"0000000111000000000000000000000000000000000000000000110000000", 		--7
	"0000111000000000000000000000000000000000000000001111000000000", 		--8
	"0000100000000000000000000000000000000000000000001000000000000", 		--9
	"0000100000000000000000000000000000000000000000001000000000000", 		--10
	"0000100000000000000000000000000000000000000000001000000000000", 		--11
	"0000100000000000000000000000000000000000000000011000000000000", 		--12
	"0000111111000000000000000000000000000000000000010000000000000", 		--13
	"0000000000100000000000000000000000000000000000011110000000000", 		--14
	"0000000000010000000000000000000000000000000000000001100000000", 		--15
	"0000000000001000000000000000000000000000000000000000010000000", 		--16
	"0000000000001000000000000000000000000000000000000000001000000",	 	--17 
	"0000000000001000000000000000000000000000000000000000000100000",		--18
	"0000000000011000000000000000000000000000000000000000000010000",		--19
	"0000000001100000000000000000000000011111111111111111111110000",		--20
	"0000000001111111111111111111111111111000000000000000000000000",		--21
	"0000000000000000000000000000000000000000000000000000000000000",		--22
	"0000000000000000000000000000000000000000000000000000000000000",		--23
	"0000000000000000000000000000000000000000000000000000000000000"		--24
	);
begin
process(rom_addra)
variable j: integer;
	begin
	     j := conv_integer(rom_addra);
   		 D <= rom(j);
end process;
end prom2_asteroid;