 library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity prom1_asteroid is
    port ( 
		rom_addra  : in std_logic_vector(7 downto 0);
        D: out STD_LOGIC_VECTOR (0 to 60)
    );
end prom1_asteroid;

architecture prom1_asteroid of prom1_asteroid is   
type rom_array is array (NATURAL range <>) of STD_LOGIC_VECTOR (0 to 60);
constant rom: rom_array := (
	"0000000000000001111111111111111111111111111110000000000000000",		--0
	"0000000000000011000000000000000000000000000001100000000000000",		--1
	"0000000000001100000000000000000000000000000001100000000000000", 		--2
	"0000000000110000000000000000000000000000000000110000000000000", 		--3
	"0000000011000000000000000000000000000000000000011000000000000", 		--4
	"0000001100000000000000000000000000000000000001100000000000000", 		--5
	"0000110000000000000000000000000000000000000001100000000000000", 		--6
	"0011000000000000000000000000000000000000000001100000000000000", 		--7
	"1100000000000000000000000000000000000000000001100000000000000", 		--8
	"1100000000000000000000000000000000000000000001100000000000000", 		--9
	"1100000000000000000000000000000000000000000000110000000000000", 		--10
	"1100000000000000000000000000000000000000000000011000000000000", 		--11
	"1100000000000000000000000000000000000000000000001100000000000", 		--12
	"0011000000000000000000000000000000000000000000000110000000000", 		--13
	"0000110000000000000000000000000000000000000000000011000000000", 		--14
	"0000001100000000000000000000000000000000000000000001100000000", 		--15
	"0000000011000000000000000000000000000000000000000001110000000", 		--16
	"0000000000110000000000000000000000000000000000000110000000000",	 	--17 
	"0000000000001100000000000000000000000000000000011000000000000",		--18
	"0000000000000011000000000000000000000000000001100000000000000",		--19
	"0000000000000000110000000000000000000000000110000000000000000",		--20
	"0000000000000000001100000000000000000000011000000000000000000",		--21
	"0000000000000000000001100000000000000001100000000000000000000",		--22
	"0000000000000000000000011111111111111110000000000000000000000",		--23
	"0000000000000000000000000000000000000000000000000000000000000"		--24
	);
begin
process(rom_addra)
variable j: integer;
	begin
	     j := conv_integer(rom_addra);
   		 D <= rom(j);
end process;
end prom1_asteroid;